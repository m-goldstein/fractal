/* This module computes the product of two complex-valued quantities by exploiting the identity that 
* (a+bi)(c+di) = (ac-bd) + i(ad+bc). Each term is computed seperately by an FPU module and then the
 * terms grouped together by ( ) are summed using another FPU module. The results from these modules 
 * is assigned to be the output values for re_z and im_z, respectively.
 */

 `include "Magic_Numbers.sv"
`define GOTO(x)				next_state = (x)

module multiplier_unit(
	input clk,
	input reset,
	input start,
	input ack,
	input [63:0] re_a,
	input [63:0] im_a,
	input [63:0] re_b,
	input [63:0] im_b,
	output logic done,
	output wire[63:0] re_z,
	output wire[63:0] im_z
	);
	
	// internal registers
	logic [63:0] ac;				// ac term (real-component of a * real-component of b)
	logic [63:0] bd;				// bd term (imaginary-component of a * imaginary-component of b)
	logic [63:0] ad;				// ad term (real-component of a * imaginary-component of b)
	logic [63:0] bc;				// bc term (imaginary-component of a * real-component of b)
	
	// internal registers for intermediate results 
	logic [63:0] _ac;
	logic [63:0] _bd;
	logic [63:0] _ad;
	logic [63:0] _bc;
	
	// logical connections (wires) to FPU modules on datapath 
	wire [63:0] re_z_wire;
	wire [63:0] im_z_wire;
	wire [63:0] ac_wire;
	wire [63:0] bd_wire;
	wire [63:0] ad_wire;
	wire [63:0] bc_wire;
	
	// internal registers for intermediate output values
	logic [63:0] re_z_out;
	logic [63:0] im_z_out;
	logic [63:0] _re_z;
	logic [63:0] _im_z;
	
	
	/* control signals */
	logic calc_re;
	logic calc_im;
	logic calc_ac;
	logic calc_bd;
	logic calc_ad;
	logic calc_bc;
	logic get_ac;
	logic get_bd; 
	logic get_ad;
	logic get_bc;
	
	logic calc_add_re;
	logic calc_add_im;	
	
	/* connections (wires) between modules on datapath */
	wire done_ac;
	wire done_bd;
	wire done_ad;
	wire done_bc;
	wire done_add_re;
	wire done_add_im;
	
	/* datapath of multiplier unit for complex values */
	/* signals to control flow of data and results within/between modules generated by control unit. */
	
	
	// define logical connections between internal registers and intermediate values of computations;
	assign ac = _ac;
	assign bd = _bd;
	assign ad = _ad;
	assign bc = _bc;
	assign re_z = re_z_out;
	assign im_z = im_z_out;
	
	// compute ac-term
	double_multiplier ac_term (
						.clk(clk),
						.reset(reset),
						.a_in(re_a),
						.b_in(re_b),
						.a_in_done(calc_ac),
						.b_in_done(calc_ac),
						.z_out_done(done_ac),
						.z_out_ack(get_ac),
						.z_out(ac_wire)
						);
						
	// compute bd-term 					
	double_multiplier bd_term (
						.clk(clk),
						.reset(reset),
						.a_in(im_a),
						.b_in(im_b),
						.a_in_done(calc_bd),
						.b_in_done(calc_bd),
						.z_out_done(done_bd),
						.z_out_ack(get_bd),
						.z_out(bd_wire)
						);
	
	// compute ad-term
	double_multiplier ad_term (
						.clk(clk),
						.reset(reset),
						.a_in(re_a),
						.b_in(im_b),
						.a_in_done(calc_ad),
						.b_in_done(calc_ad),
						.z_out_done(done_ad),
						.z_out_ack(get_ad),
						.z_out(ad_wire)
						);
						
	// compute bc-term					
	double_multiplier bc_term (
						.clk(clk),
						.reset(reset),
						.a_in(im_a),
						.b_in(re_b),
						.a_in_done(calc_bc),
						.b_in_done(calc_bc),
						.z_out_done(done_bc),
						.z_out_ack(get_bc),
						.z_out(bc_wire)
						);
						
	// compute real-component by summing ac- and bd-terms.					
	double_adder re_sum (
					.clk(clk),
					.reset(reset),
					.a_in(_ac),
					.b_in(_bd | `NEG_BITMASK),
					.a_in_done(calc_add_re),
					.b_in_done(calc_add_re),
					.z_out_ack(calc_re),
					.z_out(re_z_wire),
					.z_out_done(done_add_re)
					);
	
	// compute imaginary-component by summing ad- and bc-terms.
	double_adder im_sum (
					.clk(clk),
					.reset(reset),
					.a_in(_ad),
					.b_in(_bc),
					.a_in_done(calc_add_im),
					.b_in_done(calc_add_im),
					.z_out_ack(calc_im),
					.z_out(im_z_wire),
					.z_out_done(done_add_im)
					);
					
	enum logic[3:0] {
		HALT,
		COMPUTE_CROSS_TERMS,
		ACK_CROSS_TERMS,
		COMPUTE_COMPLEX_COMPONENTS,
		ACK_COMPLEX_COMPONENTS
	} state, next_state;
	
	always_ff @ (posedge clk) begin
		state <= (reset) ? HALT : next_state;
		_re_z <= (reset) ? `ZERO : re_z_out;
		_im_z <= (reset) ? `ZERO : im_z_out;
	end
	
	/* control logic progresses through steps of term-by-term computation of complex-valued product. */
	/* first, terms representing ac, bd, ad, bc, are computed. then real- and imaginary components are summed to form the result. */
	always_comb begin
	next_state = state;
	
	// default control signal values
	calc_add_re = 0;
	calc_add_im = 0;
	calc_ac = 0;
	calc_bd = 0;
	calc_ad = 0;
	calc_bc = 0;
	get_ac = 0;
	get_bd = 0;
	get_ad = 0;
	get_bc = 0;
	calc_re = 0;
	calc_im = 0;
	done = 0;
	
	// default assignments
	_ac = ac;
	_bd = bd;
	_ad = ad;
	_bc = bc;
	re_z_out = _re_z;
	im_z_out = _im_z;
	
	case (state)
		HALT: begin
			_ac = `ZERO;
			_bd = `ZERO;
			_ad = `ZERO;
			_bc = `ZERO;
			re_z_out = `ZERO;
			im_z_out = `ZERO;
			`GOTO( (start) ? COMPUTE_CROSS_TERMS : HALT);						// wait for start signal from generate_fractal module.
		end
		
		COMPUTE_CROSS_TERMS: begin
			// invoke multiplier units to perform computations for terms
			calc_ac = 1;
			calc_bd = 1;
			calc_ad = 1;
			calc_bc = 1;
			`GOTO ( (done_ac && done_bd && done_ad && done_bc) ? ACK_CROSS_TERMS : COMPUTE_CROSS_TERMS); // stall until all terms are computed by FPU modules.
		end
		
		ACK_CROSS_TERMS: begin
			// send ack signals to multiplier units
			get_ac = 1;
			get_bd = 1;
			get_ad = 1;
			get_bc = 1;
			
			// load outputs from ac-,bd-,ad-,bc-term modules into internal registers for intermediate processing
			_ac = ac_wire;
			_bd = bd_wire;
			_ad = ad_wire;
			_bc = bc_wire;
			`GOTO (COMPUTE_COMPLEX_COMPONENTS);						// proceed to next step and sum each complex component.
		end
		
		COMPUTE_COMPLEX_COMPONENTS: begin
			// invoke adder units to sum complex-components.
			calc_add_re = 1;
			calc_add_im = 1;
			`GOTO( (done_add_re && done_add_im) ? ACK_COMPLEX_COMPONENTS : COMPUTE_COMPLEX_COMPONENTS);	// stall until sums of both components are computed
			
		end
		
		ACK_COMPLEX_COMPONENTS: begin
			// send ack/done signals to adder units and upper-level datapath.
			calc_re = 1;
			calc_im = 1;
			done = 1;
			
			// load adder unit outputs into internal registers for intermediate result processing.
			re_z_out = re_z_wire;
			im_z_out = im_z_wire;
			`GOTO ( (ack) ? HALT : ACK_COMPLEX_COMPONENTS);				// wait for next rising edge of acknowledgement to begin next computation cycle.
			
		end
	endcase
end
endmodule
